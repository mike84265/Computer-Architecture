module Hazard_Detection (
    ID_EX_MemRd_i, ID_EX_Rt_i,
    IF_ID_Rs_i, IF_ID_Rt_i,
    Stall_o
);
